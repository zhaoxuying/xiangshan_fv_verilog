//commit 4a699e275a42daaf03e4f014bad0bb16d893e6ff
//Author: zhanglinjuan <zhanglinjuan16@mails.ucas.ac.cn>
//Date:   Tue Feb 25 10:23:28 2025 +0800
//
//    feat: support seperate DebugModule TileLink bus (#4299)
//    
//    This commit supports a configurable extra TileLink bus for DebugModule
//    besides the peripheral device bus. This involves all 3 environments
//    including TileLink-XSTop, CHI-XSTop, CHI-XSNoCTop. The feature is
//    disabled by default. To enable it, you can add `SEPERATE_DM_BUS=1` in
//    the make command line.
// Generated by CIRCT firtool-1.62.1
// Standard header to adapt well known macros for register randomization.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module SimTop(
  input         clock,
  input         reset,
  output [63:0] difftest_exit,
  output [63:0] difftest_step,
  input         difftest_perfCtrl_clean,
  input         difftest_perfCtrl_dump,
  input  [63:0] difftest_logCtrl_begin,
  input  [63:0] difftest_logCtrl_end,
  input  [63:0] difftest_logCtrl_level,
  output        difftest_uart_out_valid,
  output [7:0]  difftest_uart_out_ch,
  output        difftest_uart_in_valid,
  input  [7:0]  difftest_uart_in_ch
);


assign difftest_uart_out_valid = 0;
assign difftest_uart_out_ch = 0;
assign difftest_uart_in_valid = 0;


assign difftest_exit = 64'h0;
assign difftest_step = 64'h1;

wire  r_enable;
wire [63:0] r_index;
wire [63:0] r_data_0;
wire [63:0] r_data_1;
wire [63:0] r_data_2;
wire [63:0] r_data_3;
wire         _difftest_delayer_o_valid  ;
wire         _difftest_delayer_1_o_valid;
wire         _difftest_delayer_2_o_valid;
wire         _difftest_delayer_3_o_valid;
wire         _difftest_delayer_4_o_valid;
wire         _difftest_delayer_5_o_valid;
wire         _difftest_delayer_6_o_valid;
wire         _difftest_delayer_7_o_valid;
wire         _difftest_delayer_o_rfwen  ;
wire         _difftest_delayer_1_o_rfwen;
wire         _difftest_delayer_2_o_rfwen;
wire         _difftest_delayer_3_o_rfwen;
wire         _difftest_delayer_4_o_rfwen;
wire         _difftest_delayer_5_o_rfwen;
wire         _difftest_delayer_6_o_rfwen;
wire         _difftest_delayer_7_o_rfwen;
wire [7:0]   _difftest_delayer_o_wdest  ;
wire [7:0]   _difftest_delayer_1_o_wdest;
wire [7:0]   _difftest_delayer_2_o_wdest;
wire [7:0]   _difftest_delayer_3_o_wdest;
wire [7:0]   _difftest_delayer_4_o_wdest;
wire [7:0]   _difftest_delayer_5_o_wdest;
wire [7:0]   _difftest_delayer_6_o_wdest;
wire [7:0]   _difftest_delayer_7_o_wdest;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_0 ;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_1 ;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_2 ;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_3 ;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_4 ;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_5 ;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_6 ;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_7 ;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_8 ;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_9 ;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_10;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_11;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_12;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_13;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_14;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_15;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_16;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_17;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_18;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_19;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_20;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_21;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_22;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_23;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_24;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_25;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_26;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_27;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_28;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_29;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_30;
wire [63:0]  _difftestArchIntRegState_delayer_o_value_31;

wire commit_valid [0:7];
wire intrf_wen [0:7]; //high valid
wire [4:0] intrf_dest [0:7];
wire [63:0] intrf [0:31];

DutTop dut_top(
  .clock(clock),
  .reset(reset),
  .r_enable(r_enable),
  .r_index(r_index),
  .r_data_0(r_data_0),
  .r_data_1(r_data_1),
  .r_data_2(r_data_2),
  .r_data_3(r_data_3),
  ._difftest_delayer_o_valid  (_difftest_delayer_o_valid  ),
  ._difftest_delayer_1_o_valid(_difftest_delayer_1_o_valid),
  ._difftest_delayer_2_o_valid(_difftest_delayer_2_o_valid),
  ._difftest_delayer_3_o_valid(_difftest_delayer_3_o_valid),
  ._difftest_delayer_4_o_valid(_difftest_delayer_4_o_valid),
  ._difftest_delayer_5_o_valid(_difftest_delayer_5_o_valid),
  ._difftest_delayer_6_o_valid(_difftest_delayer_6_o_valid),
  ._difftest_delayer_7_o_valid(_difftest_delayer_7_o_valid),
  ._difftest_delayer_o_rfwen  (_difftest_delayer_o_rfwen  ),
  ._difftest_delayer_1_o_rfwen(_difftest_delayer_1_o_rfwen),
  ._difftest_delayer_2_o_rfwen(_difftest_delayer_2_o_rfwen),
  ._difftest_delayer_3_o_rfwen(_difftest_delayer_3_o_rfwen),
  ._difftest_delayer_4_o_rfwen(_difftest_delayer_4_o_rfwen),
  ._difftest_delayer_5_o_rfwen(_difftest_delayer_5_o_rfwen),
  ._difftest_delayer_6_o_rfwen(_difftest_delayer_6_o_rfwen),
  ._difftest_delayer_7_o_rfwen(_difftest_delayer_7_o_rfwen),
  ._difftest_delayer_o_wdest  (_difftest_delayer_o_wdest  ),
  ._difftest_delayer_1_o_wdest(_difftest_delayer_1_o_wdest),
  ._difftest_delayer_2_o_wdest(_difftest_delayer_2_o_wdest),
  ._difftest_delayer_3_o_wdest(_difftest_delayer_3_o_wdest),
  ._difftest_delayer_4_o_wdest(_difftest_delayer_4_o_wdest),
  ._difftest_delayer_5_o_wdest(_difftest_delayer_5_o_wdest),
  ._difftest_delayer_6_o_wdest(_difftest_delayer_6_o_wdest),
  ._difftest_delayer_7_o_wdest(_difftest_delayer_7_o_wdest),
  ._difftestArchIntRegState_delayer_o_value_0 (_difftestArchIntRegState_delayer_o_value_0 ),
  ._difftestArchIntRegState_delayer_o_value_1 (_difftestArchIntRegState_delayer_o_value_1 ),
  ._difftestArchIntRegState_delayer_o_value_2 (_difftestArchIntRegState_delayer_o_value_2 ),
  ._difftestArchIntRegState_delayer_o_value_3 (_difftestArchIntRegState_delayer_o_value_3 ),
  ._difftestArchIntRegState_delayer_o_value_4 (_difftestArchIntRegState_delayer_o_value_4 ),
  ._difftestArchIntRegState_delayer_o_value_5 (_difftestArchIntRegState_delayer_o_value_5 ),
  ._difftestArchIntRegState_delayer_o_value_6 (_difftestArchIntRegState_delayer_o_value_6 ),
  ._difftestArchIntRegState_delayer_o_value_7 (_difftestArchIntRegState_delayer_o_value_7 ),
  ._difftestArchIntRegState_delayer_o_value_8 (_difftestArchIntRegState_delayer_o_value_8 ),
  ._difftestArchIntRegState_delayer_o_value_9 (_difftestArchIntRegState_delayer_o_value_9 ),
  ._difftestArchIntRegState_delayer_o_value_10(_difftestArchIntRegState_delayer_o_value_10),
  ._difftestArchIntRegState_delayer_o_value_11(_difftestArchIntRegState_delayer_o_value_11),
  ._difftestArchIntRegState_delayer_o_value_12(_difftestArchIntRegState_delayer_o_value_12),
  ._difftestArchIntRegState_delayer_o_value_13(_difftestArchIntRegState_delayer_o_value_13),
  ._difftestArchIntRegState_delayer_o_value_14(_difftestArchIntRegState_delayer_o_value_14),
  ._difftestArchIntRegState_delayer_o_value_15(_difftestArchIntRegState_delayer_o_value_15),
  ._difftestArchIntRegState_delayer_o_value_16(_difftestArchIntRegState_delayer_o_value_16),
  ._difftestArchIntRegState_delayer_o_value_17(_difftestArchIntRegState_delayer_o_value_17),
  ._difftestArchIntRegState_delayer_o_value_18(_difftestArchIntRegState_delayer_o_value_18),
  ._difftestArchIntRegState_delayer_o_value_19(_difftestArchIntRegState_delayer_o_value_19),
  ._difftestArchIntRegState_delayer_o_value_20(_difftestArchIntRegState_delayer_o_value_20),
  ._difftestArchIntRegState_delayer_o_value_21(_difftestArchIntRegState_delayer_o_value_21),
  ._difftestArchIntRegState_delayer_o_value_22(_difftestArchIntRegState_delayer_o_value_22),
  ._difftestArchIntRegState_delayer_o_value_23(_difftestArchIntRegState_delayer_o_value_23),
  ._difftestArchIntRegState_delayer_o_value_24(_difftestArchIntRegState_delayer_o_value_24),
  ._difftestArchIntRegState_delayer_o_value_25(_difftestArchIntRegState_delayer_o_value_25),
  ._difftestArchIntRegState_delayer_o_value_26(_difftestArchIntRegState_delayer_o_value_26),
  ._difftestArchIntRegState_delayer_o_value_27(_difftestArchIntRegState_delayer_o_value_27),
  ._difftestArchIntRegState_delayer_o_value_28(_difftestArchIntRegState_delayer_o_value_28),
  ._difftestArchIntRegState_delayer_o_value_29(_difftestArchIntRegState_delayer_o_value_29),
  ._difftestArchIntRegState_delayer_o_value_30(_difftestArchIntRegState_delayer_o_value_30),
  ._difftestArchIntRegState_delayer_o_value_31(_difftestArchIntRegState_delayer_o_value_31)
);

  DifftestMem1P rdata_mem (
    .clock        (clock),
    .reset        (reset),
    .read_valid   (r_enable),
    .read_index   (r_index),
    .read_data_0  (r_data_0),
    .read_data_1  (r_data_1),
    .read_data_2  (r_data_2),
    .read_data_3  (r_data_3),
    .write_valid  (1'b0),
    .write_index  (64'b0),
    .write_data_0 (64'b0),
    .write_data_1 (64'b0),
    .write_data_2 (64'b0),
    .write_data_3 (64'b0),
    .write_mask_0 (64'b0),
    .write_mask_1 (64'b0),
    .write_mask_2 (64'b0),
    .write_mask_3 (64'b0)
  );

`ifdef TRY_DEBUG
assign commit_valid[0] = _difftest_delayer_o_valid;
assign commit_valid[1] = _difftest_delayer_1_o_valid;
assign commit_valid[2] = _difftest_delayer_2_o_valid;
assign commit_valid[3] = _difftest_delayer_3_o_valid;
assign commit_valid[4] = _difftest_delayer_4_o_valid;
assign commit_valid[5] = _difftest_delayer_5_o_valid;
assign commit_valid[6] = _difftest_delayer_6_o_valid;
assign commit_valid[7] = _difftest_delayer_7_o_valid;

assign intrf_wen[0] = _difftest_delayer_o_rfwen;
assign intrf_wen[1] = _difftest_delayer_1_o_rfwen;
assign intrf_wen[2] = _difftest_delayer_2_o_rfwen;
assign intrf_wen[3] = _difftest_delayer_3_o_rfwen;
assign intrf_wen[4] = _difftest_delayer_4_o_rfwen;
assign intrf_wen[5] = _difftest_delayer_5_o_rfwen;
assign intrf_wen[6] = _difftest_delayer_6_o_rfwen;
assign intrf_wen[7] = _difftest_delayer_7_o_rfwen;

assign intrf_dest[0] = _difftest_delayer_o_wdest[4:0];
assign intrf_dest[1] = _difftest_delayer_1_o_wdest[4:0];
assign intrf_dest[2] = _difftest_delayer_2_o_wdest[4:0];
assign intrf_dest[3] = _difftest_delayer_3_o_wdest[4:0];
assign intrf_dest[4] = _difftest_delayer_4_o_wdest[4:0];
assign intrf_dest[5] = _difftest_delayer_5_o_wdest[4:0];
assign intrf_dest[6] = _difftest_delayer_6_o_wdest[4:0];
assign intrf_dest[7] = _difftest_delayer_7_o_wdest[4:0];

assign intrf[0 ] = _difftestArchIntRegState_delayer_o_value_0 ; 
assign intrf[1 ] = _difftestArchIntRegState_delayer_o_value_1 ; 
assign intrf[2 ] = _difftestArchIntRegState_delayer_o_value_2 ; 
assign intrf[3 ] = _difftestArchIntRegState_delayer_o_value_3 ; 
assign intrf[4 ] = _difftestArchIntRegState_delayer_o_value_4 ; 
assign intrf[5 ] = _difftestArchIntRegState_delayer_o_value_5 ; 
assign intrf[6 ] = _difftestArchIntRegState_delayer_o_value_6 ; 
assign intrf[7 ] = _difftestArchIntRegState_delayer_o_value_7 ; 
assign intrf[8 ] = _difftestArchIntRegState_delayer_o_value_8 ; 
assign intrf[9 ] = _difftestArchIntRegState_delayer_o_value_9 ; 
assign intrf[10] = _difftestArchIntRegState_delayer_o_value_10; 
assign intrf[11] = _difftestArchIntRegState_delayer_o_value_11; 
assign intrf[12] = _difftestArchIntRegState_delayer_o_value_12; 
assign intrf[13] = _difftestArchIntRegState_delayer_o_value_13; 
assign intrf[14] = _difftestArchIntRegState_delayer_o_value_14; 
assign intrf[15] = _difftestArchIntRegState_delayer_o_value_15; 
assign intrf[16] = _difftestArchIntRegState_delayer_o_value_16; 
assign intrf[17] = _difftestArchIntRegState_delayer_o_value_17; 
assign intrf[18] = _difftestArchIntRegState_delayer_o_value_18; 
assign intrf[19] = _difftestArchIntRegState_delayer_o_value_19; 
assign intrf[20] = _difftestArchIntRegState_delayer_o_value_20; 
assign intrf[21] = _difftestArchIntRegState_delayer_o_value_21; 
assign intrf[22] = _difftestArchIntRegState_delayer_o_value_22; 
assign intrf[23] = _difftestArchIntRegState_delayer_o_value_23; 
assign intrf[24] = _difftestArchIntRegState_delayer_o_value_24; 
assign intrf[25] = _difftestArchIntRegState_delayer_o_value_25; 
assign intrf[26] = _difftestArchIntRegState_delayer_o_value_26; 
assign intrf[27] = _difftestArchIntRegState_delayer_o_value_27; 
assign intrf[28] = _difftestArchIntRegState_delayer_o_value_28; 
assign intrf[29] = _difftestArchIntRegState_delayer_o_value_29; 
assign intrf[30] = _difftestArchIntRegState_delayer_o_value_30; 
assign intrf[31] = _difftestArchIntRegState_delayer_o_value_31;

// EDIT: Insert the qed ready logic -- tracks number of committed instructions
(* keep *)
wire qed_ready;
(* keep *)
reg [15:0] num_orig_insts;
(* keep *)
reg [15:0] num_dup_insts;
reg [3:0] num_orig_commits;
reg [3:0] num_dup_commits;

integer fp;

initial begin
  fp = $fopen("try_debug.log", "w");
  if (fp == 0) begin
    $display("can't open try_debug.log!");
    $finish;
  end
end

always @(*) begin
  num_orig_commits = 0;
  for (int i = 0; i < 8; i = i + 1) begin
    if (commit_valid[i] && intrf_wen[i] && (intrf_dest[i] < 5'd16) && (intrf_dest[i] != 0))
      num_orig_commits = num_orig_commits + 1;
  end
end

always @(*) begin
  num_dup_commits = 0;
  for (int i = 0; i < 8; i = i + 1) begin
    if (commit_valid[i] && intrf_wen[i] && (intrf_dest[i] >= 5'd16))
      num_dup_commits = num_dup_commits + 1;
  end
end

always @(posedge clock) begin
  if (reset) begin
    num_orig_insts <= 16'b0;
    num_dup_insts <= 16'b0;
  end 
  else begin
    num_orig_insts <= num_orig_insts + {12'b0,num_orig_commits};
    num_dup_insts <= num_dup_insts + {12'b0,num_dup_commits};
  end
end

assign qed_ready = (num_orig_insts == num_dup_insts);

always @(posedge clock) begin
  if(num_orig_insts!=16'b0 || num_dup_insts!=16'b0) begin
    $fdisplay(fp, "num_orig_commits = %6d, num_orig_insts = %6d,      num_dup_commits = %6d, num_dup_insts = %6d",num_orig_commits,num_orig_insts,num_dup_commits,num_dup_insts);
    $fdisplay(fp, "intrf1=%016h, intrf17=%016h",intrf[1],intrf[17]);
  end
end

final begin
  $fclose(fp);
end
`endif //TRY_DEBUG

endmodule

